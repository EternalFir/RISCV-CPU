`include "constants.v"
`include "Decoder.v"

module Dispatcher(

);

endmodule : Dispatcher